package or_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    import seq_item_pkg::*;
    `include "or_agent_config.svh"
    `include "or_sequencer.svh"
    `include "or_driver.svh"
    `include "or_monitor.svh"
    `include "or_agent.svh"
        
endpackage :or_agent_pkg