package v_seq_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    `include "virtual_sequence.svh"
    `include "v_random_seq.svh"
    `include "v_all_zero_seq.svh"
    `include "v_all_one_seq.svh"
endpackage :v_seq_pkg