package and_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    import seq_item_pkg::*;
    `include "and_agent_config.svh"
    `include "and_sequencer.svh"
    `include "and_driver.svh"
    `include "and_monitor.svh"
    `include "and_agent.svh"
        
endpackage :and_agent_pkg