package seq_item_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;
    `include "and_seq_item.svh"
    `include "or_seq_item.svh"
    `include "shift_seq_item.svh"
    `include "xor_seq_item.svh"
    
endpackage :seq_item_pkg