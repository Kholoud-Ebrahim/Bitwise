class or_all_one_seq extends or_base_seq;
    `uvm_object_utils(or_all_one_seq)

    or_seq_item  or_item;

    function new(string name = "or_all_one_seq");
        super.new(name);
    endfunction

    task body();
        or_item = or_seq_item::type_id::create("or_item");
        start_item(or_item);
        assert(or_item.randomize() with {or_in1 == {OWIDTH{1'b1}}; or_in2 == {OWIDTH{1'b1}};});
        finish_item(or_item);
    endtask :body
endclass :or_all_one_seq