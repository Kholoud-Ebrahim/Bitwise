package test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import param_pkg::*;

    `include "base_test.svh"
    `include "random_test.svh"
    `include "all_zero_test.svh"
    `include "all_one_test.svh"
endpackage :test_pkg