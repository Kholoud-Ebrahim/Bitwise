package param_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    parameter PERIOD = 20;
    parameter AWIDTH =8;
    parameter OWIDTH =8;
    parameter XWIDTH =8;
    parameter SRWIDTH =8, SROPWIDTH =8;
    parameter SLWIDTH =8, SLOPWIDTH =8;
endpackage :param_pkg